library ieee;
use ieee.std_logic_1164.ALL;

package definitions is
	type t_pattern is (no_pattern, first_one, second_zero, second_one, pattern_rec);
end definitions;

package body definitions is

end definitions;
